module Final_Project_287(clk, rst);
	
	
	
endmodule 